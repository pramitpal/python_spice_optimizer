***** 2nd Order RC Circuit Frequency Response *****
.PARAM R_1 = 1200.0
.PARAM C_1 = 1e-06
.PARAM START = 1
.PARAM STOP = 1000000000.0
**--**--**--**--**--**--**--**--**--**
r1 1 2 {R_1}
c1 2 0 {C_1}


********Specifying an AC source with zero dc
vin 1 0 dc 0 ac 1
********AC analysis for 1 Hz to 1MHz, 10 points per decade
.ac dec 10 {START} {STOP}


.control
set filetype=ascii
run

let m=vdb(2)

*plot m xlog

meas ac cutoff find frequency WHEN m=-3.0 CROSS=LAST

write rc_test.raw cutoff
.endc
.end
